<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>8.65382,0.484882,83.6632,-37.8636</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>31,-21</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>31,-30</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>31,-25</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>29,-21</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>29,-24.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>29,-29.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>31,-7</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>31,-9</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>31,-14</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>37,-22</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_AND2</type>
<position>37,-27</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_OR3</type>
<position>46.5,-27</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>30 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>69</ID>
<type>GA_LED</type>
<position>52,-27</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>29,-6.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>29,-9</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>29,-14</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>37,-8</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR2</type>
<position>43,-10.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>52,-10.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>48,-17</position>
<gparam>LABEL_TEXT -------------------------------------------------------------------------------------</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-26,34,-23</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,-25,34,-25</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>33,-21,34,-21</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>34 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>34,-21,34,-21</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-21 4</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-30,43.5,-30</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>34 6</intersection>
<intersection>43.5 10</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>34,-30,34,-28</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>43.5,-30,43.5,-29</points>
<connection>
<GID>67</GID>
<name>IN_2</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-25,40,-22</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>40,-25,43.5,-25</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-27,43.5,-27</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-27,51,-27</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>33,-7,34,-7</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-9,34,-9</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-9.5,40,-8</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-14,36.5,-11.5</points>
<intersection>-14 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-11.5,40,-11.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-14,36.5,-14</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-10.5,51,-10.5</points>
<connection>
<GID>78</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 9></circuit>